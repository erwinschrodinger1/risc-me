module main();

initial
  begin
    
  end

endmodule